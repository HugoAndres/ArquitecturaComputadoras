// PLL.v

// Generated using ACDS version 12.1 177 at 2021.12.14.23:11:32

`timescale 1 ps / 1 ps
module PLL (
		input  wire  clkin_clk,   //   clkin.clk
		output wire  clkout2_clk, // clkout2.clk
		input  wire  reset_reset, //   reset.reset
		output wire  clkout1_clk  // clkout1.clk
	);

	PLL_altpll_0 altpll_0 (
		.clk       (clkin_clk),   //       inclk_interface.clk
		.reset     (reset_reset), // inclk_interface_reset.reset
		.read      (),            //             pll_slave.read
		.write     (),            //                      .write
		.address   (),            //                      .address
		.readdata  (),            //                      .readdata
		.writedata (),            //                      .writedata
		.c0        (clkout1_clk), //                    c0.clk
		.c1        (clkout2_clk), //                    c1.clk
		.areset    (),            //        areset_conduit.export
		.locked    (),            //        locked_conduit.export
		.phasedone ()             //     phasedone_conduit.export
	);

endmodule
